module por_rosc (clk_8mhz,
    clk_out,
    fb_in,
    fb_out,
    one,
    por_n,
    rst_n,
    zero,
    VGND,
    VPWR,
    freq_sel);
 output clk_8mhz;
 output clk_out;
 input fb_in;
 output fb_out;
 input one;
 output por_n;
 input rst_n;
 input zero;
 input VGND;
 input VPWR;
 input [1:0] freq_sel;

 wire \CLKMUX.clk1 ;
 wire \CLKMUX.clk2 ;
 wire \CLKMUX.clk3 ;
 wire \CLKMUX.clk4 ;
 wire \CLKMUX.m1.Q1a ;
 wire \CLKMUX.m1.Q1b ;
 wire \CLKMUX.m1.Q2a ;
 wire \CLKMUX.m1.Q2b ;
 wire \CLKMUX.m1.q1a_in ;
 wire \CLKMUX.m1.q2a_in ;
 wire \CLKMUX.m2.Q1a ;
 wire \CLKMUX.m2.Q1b ;
 wire \CLKMUX.m2.Q2a ;
 wire \CLKMUX.m2.Q2b ;
 wire \CLKMUX.m2.q1a_in ;
 wire \CLKMUX.m2.q2a_in ;
 wire \CLKMUX.m3.Q1a ;
 wire \CLKMUX.m3.Q1b ;
 wire \CLKMUX.m3.Q2a ;
 wire \CLKMUX.m3.Q2b ;
 wire \CLKMUX.m3.q1a_in ;
 wire \CLKMUX.m3.q2a_in ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire \clk_div[1] ;
 wire \clk_div[2] ;
 wire \clk_div[3] ;
 wire \clk_div[4] ;
 wire \clk_div[5] ;
 wire \clk_div[6] ;
 wire \clk_div[7] ;
 wire \clk_div[8] ;
 wire cmp0;
 wire cmp1;
 wire cmp2;
 wire cmp3;
 wire \dly[1] ;
 wire \dly[2] ;
 wire \dly[3] ;
 wire \dly[4] ;
 wire \dly[5] ;
 wire \dly[6] ;
 wire \dly[7] ;
 wire \shift_reg0[0] ;
 wire \shift_reg0[10] ;
 wire \shift_reg0[11] ;
 wire \shift_reg0[12] ;
 wire \shift_reg0[13] ;
 wire \shift_reg0[14] ;
 wire \shift_reg0[15] ;
 wire \shift_reg0[1] ;
 wire \shift_reg0[2] ;
 wire \shift_reg0[3] ;
 wire \shift_reg0[4] ;
 wire \shift_reg0[5] ;
 wire \shift_reg0[6] ;
 wire \shift_reg0[7] ;
 wire \shift_reg0[8] ;
 wire \shift_reg0[9] ;
 wire \shift_reg1[0] ;
 wire \shift_reg1[10] ;
 wire \shift_reg1[11] ;
 wire \shift_reg1[12] ;
 wire \shift_reg1[13] ;
 wire \shift_reg1[14] ;
 wire \shift_reg1[15] ;
 wire \shift_reg1[1] ;
 wire \shift_reg1[2] ;
 wire \shift_reg1[3] ;
 wire \shift_reg1[4] ;
 wire \shift_reg1[5] ;
 wire \shift_reg1[6] ;
 wire \shift_reg1[7] ;
 wire \shift_reg1[8] ;
 wire \shift_reg1[9] ;
 wire \shift_reg2[0] ;
 wire \shift_reg2[10] ;
 wire \shift_reg2[11] ;
 wire \shift_reg2[12] ;
 wire \shift_reg2[13] ;
 wire \shift_reg2[14] ;
 wire \shift_reg2[15] ;
 wire \shift_reg2[1] ;
 wire \shift_reg2[2] ;
 wire \shift_reg2[3] ;
 wire \shift_reg2[4] ;
 wire \shift_reg2[5] ;
 wire \shift_reg2[6] ;
 wire \shift_reg2[7] ;
 wire \shift_reg2[8] ;
 wire \shift_reg2[9] ;
 wire \shift_reg3[0] ;
 wire \shift_reg3[10] ;
 wire \shift_reg3[11] ;
 wire \shift_reg3[12] ;
 wire \shift_reg3[13] ;
 wire \shift_reg3[14] ;
 wire \shift_reg3[15] ;
 wire \shift_reg3[1] ;
 wire \shift_reg3[2] ;
 wire \shift_reg3[3] ;
 wire \shift_reg3[4] ;
 wire \shift_reg3[5] ;
 wire \shift_reg3[6] ;
 wire \shift_reg3[7] ;
 wire \shift_reg3[8] ;
 wire \shift_reg3[9] ;

 sky130_fd_sc_hs__clkbuf_8 CLKBUF_0 (.A(\dly[7] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(fb_out));
 sky130_fd_sc_hs__clkbuf_4 CLKBUF_1 (.A(fb_out),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(\CLKMUX.clk1 ));
 sky130_fd_sc_hs__clkdlyinv5sd3_1 DLYINV_0 (.A(fb_in),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\dly[1] ));
 sky130_fd_sc_hs__clkdlyinv5sd3_1 DLYINV_1 (.A(\dly[1] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\dly[2] ));
 sky130_fd_sc_hs__clkdlyinv5sd3_1 DLYINV_2 (.A(\dly[2] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\dly[3] ));
 sky130_fd_sc_hs__clkdlyinv5sd3_1 DLYINV_3 (.A(\dly[3] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\dly[4] ));
 sky130_fd_sc_hs__clkdlyinv5sd3_1 DLYINV_4 (.A(\dly[4] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\dly[5] ));
 sky130_fd_sc_hs__clkdlyinv5sd2_1 DLYINV_5 (.A(\dly[5] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\dly[6] ));
 sky130_fd_sc_hs__clkdlyinv5sd2_1 DLYINV_6 (.A(\dly[6] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\dly[7] ));
 sky130_fd_sc_hs__clkinv_1 _075_ (.A(\CLKMUX.clk2 ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_002_));
 sky130_fd_sc_hs__clkinv_1 _076_ (.A(\CLKMUX.m3.Q1b ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_010_));
 sky130_fd_sc_hs__clkinv_1 _077_ (.A(\CLKMUX.m3.Q2b ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_011_));
 sky130_fd_sc_hs__nand3_1 _078_ (.A(\shift_reg0[9] ),
    .B(\shift_reg0[10] ),
    .C(\shift_reg0[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_012_));
 sky130_fd_sc_hs__nand2_1 _079_ (.A(one),
    .B(\shift_reg0[4] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_013_));
 sky130_fd_sc_hs__nand4_1 _080_ (.A(\shift_reg0[5] ),
    .B(\shift_reg0[6] ),
    .C(\shift_reg0[7] ),
    .D(\shift_reg0[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_014_));
 sky130_fd_sc_hs__nor3_1 _081_ (.A(_012_),
    .B(_013_),
    .C(_014_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_015_));
 sky130_fd_sc_hs__nor3_1 _082_ (.A(\shift_reg0[9] ),
    .B(\shift_reg0[10] ),
    .C(\shift_reg0[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_016_));
 sky130_fd_sc_hs__or4_1 _083_ (.A(one),
    .B(\shift_reg0[4] ),
    .C(\shift_reg0[5] ),
    .D(\shift_reg0[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_017_));
 sky130_fd_sc_hs__nor4b_1 _084_ (.A(\shift_reg0[6] ),
    .B(_017_),
    .C(\shift_reg0[7] ),
    .D_N(_016_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_018_));
 sky130_fd_sc_hs__nand2_1 _085_ (.A(\shift_reg0[1] ),
    .B(one),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_019_));
 sky130_fd_sc_hs__nand3_1 _086_ (.A(\shift_reg0[2] ),
    .B(\shift_reg0[3] ),
    .C(\shift_reg0[0] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_020_));
 sky130_fd_sc_hs__or4_1 _087_ (.A(\shift_reg0[1] ),
    .B(one),
    .C(\shift_reg0[2] ),
    .D(\shift_reg0[3] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_021_));
 sky130_fd_sc_hs__o22ai_1 _088_ (.A1(_019_),
    .A2(_020_),
    .B1(_021_),
    .B2(\shift_reg0[0] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_022_));
 sky130_fd_sc_hs__nand2_1 _089_ (.A(one),
    .B(\shift_reg0[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_023_));
 sky130_fd_sc_hs__nand3_1 _090_ (.A(\shift_reg0[13] ),
    .B(\shift_reg0[14] ),
    .C(\shift_reg0[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_024_));
 sky130_fd_sc_hs__or4_1 _091_ (.A(one),
    .B(\shift_reg0[12] ),
    .C(\shift_reg0[13] ),
    .D(\shift_reg0[14] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_025_));
 sky130_fd_sc_hs__o22ai_1 _092_ (.A1(_023_),
    .A2(_024_),
    .B1(_025_),
    .B2(\shift_reg0[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_026_));
 sky130_fd_sc_hs__o211a_2 _093_ (.A1(_015_),
    .A2(_018_),
    .B1(_022_),
    .C1(_026_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(cmp0));
 sky130_fd_sc_hs__and3_1 _094_ (.A(\shift_reg1[9] ),
    .B(\shift_reg1[10] ),
    .C(\shift_reg1[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_027_));
 sky130_fd_sc_hs__and4_1 _095_ (.A(zero),
    .B(\shift_reg1[4] ),
    .C(\shift_reg1[5] ),
    .D(\shift_reg1[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_028_));
 sky130_fd_sc_hs__nand4_1 _096_ (.A(\shift_reg1[6] ),
    .B(\shift_reg1[7] ),
    .C(_027_),
    .D(_028_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_029_));
 sky130_fd_sc_hs__nor3_1 _097_ (.A(\shift_reg1[9] ),
    .B(\shift_reg1[10] ),
    .C(\shift_reg1[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_030_));
 sky130_fd_sc_hs__nor2_1 _098_ (.A(zero),
    .B(\shift_reg1[4] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_031_));
 sky130_fd_sc_hs__nor4_1 _099_ (.A(\shift_reg1[5] ),
    .B(\shift_reg1[6] ),
    .C(\shift_reg1[7] ),
    .D(\shift_reg1[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_032_));
 sky130_fd_sc_hs__nand3_1 _100_ (.A(_030_),
    .B(_031_),
    .C(_032_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_033_));
 sky130_fd_sc_hs__nor3_1 _101_ (.A(\shift_reg1[13] ),
    .B(\shift_reg1[14] ),
    .C(\shift_reg1[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_034_));
 sky130_fd_sc_hs__nor2_1 _102_ (.A(zero),
    .B(\shift_reg1[0] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_035_));
 sky130_fd_sc_hs__nor4_1 _103_ (.A(\shift_reg1[1] ),
    .B(\shift_reg1[2] ),
    .C(\shift_reg1[3] ),
    .D(\shift_reg1[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_036_));
 sky130_fd_sc_hs__nand3_1 _104_ (.A(_034_),
    .B(_035_),
    .C(_036_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_037_));
 sky130_fd_sc_hs__and3_1 _105_ (.A(\shift_reg1[13] ),
    .B(\shift_reg1[14] ),
    .C(\shift_reg1[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_038_));
 sky130_fd_sc_hs__and4_1 _106_ (.A(\shift_reg1[1] ),
    .B(\shift_reg1[2] ),
    .C(\shift_reg1[3] ),
    .D(\shift_reg1[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_039_));
 sky130_fd_sc_hs__nand4_1 _107_ (.A(zero),
    .B(\shift_reg1[0] ),
    .C(_038_),
    .D(_039_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_040_));
 sky130_fd_sc_hs__a22oi_1 _108_ (.A1(_029_),
    .A2(_033_),
    .B1(_037_),
    .B2(_040_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(cmp1));
 sky130_fd_sc_hs__and3_1 _109_ (.A(\shift_reg2[9] ),
    .B(\shift_reg2[10] ),
    .C(\shift_reg2[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_041_));
 sky130_fd_sc_hs__and4_1 _110_ (.A(one),
    .B(\shift_reg2[4] ),
    .C(\shift_reg2[5] ),
    .D(\shift_reg2[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_042_));
 sky130_fd_sc_hs__nand4_1 _111_ (.A(\shift_reg2[6] ),
    .B(\shift_reg2[7] ),
    .C(_041_),
    .D(_042_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_043_));
 sky130_fd_sc_hs__nor3_1 _112_ (.A(\shift_reg2[9] ),
    .B(\shift_reg2[10] ),
    .C(\shift_reg2[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_044_));
 sky130_fd_sc_hs__nor2_1 _113_ (.A(one),
    .B(\shift_reg2[4] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_045_));
 sky130_fd_sc_hs__nor4_1 _114_ (.A(\shift_reg2[5] ),
    .B(\shift_reg2[6] ),
    .C(\shift_reg2[7] ),
    .D(\shift_reg2[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_046_));
 sky130_fd_sc_hs__nand3_1 _115_ (.A(_044_),
    .B(_045_),
    .C(_046_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_047_));
 sky130_fd_sc_hs__nor3_1 _116_ (.A(\shift_reg2[13] ),
    .B(\shift_reg2[14] ),
    .C(\shift_reg2[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_048_));
 sky130_fd_sc_hs__nor2_1 _117_ (.A(one),
    .B(\shift_reg2[0] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_049_));
 sky130_fd_sc_hs__nor4_1 _118_ (.A(\shift_reg2[1] ),
    .B(\shift_reg2[2] ),
    .C(\shift_reg2[3] ),
    .D(\shift_reg2[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_050_));
 sky130_fd_sc_hs__nand3_1 _119_ (.A(_048_),
    .B(_049_),
    .C(_050_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_051_));
 sky130_fd_sc_hs__and3_1 _120_ (.A(\shift_reg2[13] ),
    .B(\shift_reg2[14] ),
    .C(\shift_reg2[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_052_));
 sky130_fd_sc_hs__and4_1 _121_ (.A(\shift_reg2[1] ),
    .B(\shift_reg2[2] ),
    .C(\shift_reg2[3] ),
    .D(\shift_reg2[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_053_));
 sky130_fd_sc_hs__nand4_1 _122_ (.A(one),
    .B(\shift_reg2[0] ),
    .C(_052_),
    .D(_053_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_054_));
 sky130_fd_sc_hs__a22oi_1 _123_ (.A1(_043_),
    .A2(_047_),
    .B1(_051_),
    .B2(_054_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(cmp2));
 sky130_fd_sc_hs__and3_1 _124_ (.A(\shift_reg3[9] ),
    .B(\shift_reg3[10] ),
    .C(\shift_reg3[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_055_));
 sky130_fd_sc_hs__and4_1 _125_ (.A(zero),
    .B(\shift_reg3[4] ),
    .C(\shift_reg3[5] ),
    .D(\shift_reg3[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_056_));
 sky130_fd_sc_hs__nand4_1 _126_ (.A(\shift_reg3[6] ),
    .B(\shift_reg3[7] ),
    .C(_055_),
    .D(_056_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_057_));
 sky130_fd_sc_hs__nor3_1 _127_ (.A(\shift_reg3[9] ),
    .B(\shift_reg3[10] ),
    .C(\shift_reg3[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_058_));
 sky130_fd_sc_hs__nor2_1 _128_ (.A(zero),
    .B(\shift_reg3[4] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_059_));
 sky130_fd_sc_hs__nor4_1 _129_ (.A(\shift_reg3[5] ),
    .B(\shift_reg3[6] ),
    .C(\shift_reg3[7] ),
    .D(\shift_reg3[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_060_));
 sky130_fd_sc_hs__nand3_1 _130_ (.A(_058_),
    .B(_059_),
    .C(_060_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_061_));
 sky130_fd_sc_hs__nor3_1 _131_ (.A(\shift_reg3[13] ),
    .B(\shift_reg3[14] ),
    .C(\shift_reg3[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_062_));
 sky130_fd_sc_hs__nor2_1 _132_ (.A(zero),
    .B(\shift_reg3[0] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_063_));
 sky130_fd_sc_hs__nor4_1 _133_ (.A(\shift_reg3[1] ),
    .B(\shift_reg3[2] ),
    .C(\shift_reg3[3] ),
    .D(\shift_reg3[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_064_));
 sky130_fd_sc_hs__nand3_1 _134_ (.A(_062_),
    .B(_063_),
    .C(_064_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_065_));
 sky130_fd_sc_hs__and3_1 _135_ (.A(\shift_reg3[13] ),
    .B(\shift_reg3[14] ),
    .C(\shift_reg3[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_066_));
 sky130_fd_sc_hs__and4_1 _136_ (.A(\shift_reg3[1] ),
    .B(\shift_reg3[2] ),
    .C(\shift_reg3[3] ),
    .D(\shift_reg3[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_067_));
 sky130_fd_sc_hs__nand4_1 _137_ (.A(zero),
    .B(\shift_reg3[0] ),
    .C(_066_),
    .D(_067_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_068_));
 sky130_fd_sc_hs__a22oi_1 _138_ (.A1(_057_),
    .A2(_061_),
    .B1(_065_),
    .B2(_068_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(cmp3));
 sky130_fd_sc_hs__and4_1 _139_ (.A(cmp0),
    .B(cmp1),
    .C(cmp2),
    .D(cmp3),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(por_n));
 sky130_fd_sc_hs__a22oi_1 _140_ (.A1(\CLKMUX.clk3 ),
    .A2(\CLKMUX.m2.Q1b ),
    .B1(\CLKMUX.clk4 ),
    .B2(\CLKMUX.m2.Q2b ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_000_));
 sky130_fd_sc_hs__a22oi_1 _141_ (.A1(\CLKMUX.clk1 ),
    .A2(\CLKMUX.m1.Q1b ),
    .B1(\CLKMUX.m1.Q2b ),
    .B2(\CLKMUX.clk2 ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_001_));
 sky130_fd_sc_hs__o22ai_1 _142_ (.A1(_011_),
    .A2(_000_),
    .B1(_001_),
    .B2(_010_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(clk_out));
 sky130_fd_sc_hs__nor2_1 _143_ (.A(\CLKMUX.m3.Q2b ),
    .B(freq_sel[1]),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\CLKMUX.m3.q1a_in ));
 sky130_fd_sc_hs__nor2b_1 _144_ (.A(\CLKMUX.m3.Q1b ),
    .B_N(freq_sel[1]),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\CLKMUX.m3.q2a_in ));
 sky130_fd_sc_hs__nor2_1 _145_ (.A(\CLKMUX.m2.Q2b ),
    .B(freq_sel[0]),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\CLKMUX.m2.q1a_in ));
 sky130_fd_sc_hs__nor2b_1 _146_ (.A(\CLKMUX.m2.Q1b ),
    .B_N(freq_sel[0]),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\CLKMUX.m2.q2a_in ));
 sky130_fd_sc_hs__nor2_1 _147_ (.A(\CLKMUX.m1.Q2b ),
    .B(freq_sel[0]),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\CLKMUX.m1.q1a_in ));
 sky130_fd_sc_hs__nor2b_1 _148_ (.A(\CLKMUX.m1.Q1b ),
    .B_N(freq_sel[0]),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(\CLKMUX.m1.q2a_in ));
 sky130_fd_sc_hs__nand2_1 _149_ (.A(\CLKMUX.clk2 ),
    .B(\CLKMUX.clk3 ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_069_));
 sky130_fd_sc_hs__xnor2_1 _150_ (.A(_002_),
    .B(\CLKMUX.clk3 ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_003_));
 sky130_fd_sc_hs__xnor2_1 _151_ (.A(\CLKMUX.clk4 ),
    .B(_069_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_004_));
 sky130_fd_sc_hs__and4_1 _152_ (.A(\CLKMUX.clk2 ),
    .B(\CLKMUX.clk3 ),
    .C(\CLKMUX.clk4 ),
    .D(clk_8mhz),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_070_));
 sky130_fd_sc_hs__a31oi_1 _153_ (.A1(\CLKMUX.clk2 ),
    .A2(\CLKMUX.clk3 ),
    .A3(\CLKMUX.clk4 ),
    .B1(clk_8mhz),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_071_));
 sky130_fd_sc_hs__nor2_1 _154_ (.A(_070_),
    .B(_071_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_005_));
 sky130_fd_sc_hs__nand2_1 _155_ (.A(\clk_div[5] ),
    .B(_070_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_072_));
 sky130_fd_sc_hs__xor2_1 _156_ (.A(\clk_div[5] ),
    .B(_070_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hs__nand3_1 _157_ (.A(\clk_div[5] ),
    .B(\clk_div[6] ),
    .C(_070_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_073_));
 sky130_fd_sc_hs__xnor2_1 _158_ (.A(\clk_div[6] ),
    .B(_072_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_007_));
 sky130_fd_sc_hs__nand4_1 _159_ (.A(\clk_div[5] ),
    .B(\clk_div[6] ),
    .C(\clk_div[7] ),
    .D(_070_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_074_));
 sky130_fd_sc_hs__xnor2_1 _160_ (.A(\clk_div[7] ),
    .B(_073_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_008_));
 sky130_fd_sc_hs__xnor2_1 _161_ (.A(\clk_div[8] ),
    .B(_074_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Y(_009_));
 sky130_fd_sc_hs__dfxtp_1 _162_ (.CLK(\CLKMUX.clk1 ),
    .D(_002_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.clk2 ));
 sky130_fd_sc_hs__dfxtp_1 _163_ (.CLK(\CLKMUX.clk1 ),
    .D(_003_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.clk3 ));
 sky130_fd_sc_hs__dfxtp_1 _164_ (.CLK(\CLKMUX.clk1 ),
    .D(_004_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.clk4 ));
 sky130_fd_sc_hs__dfxtp_1 _165_ (.CLK(\CLKMUX.clk1 ),
    .D(_005_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(clk_8mhz));
 sky130_fd_sc_hs__dfxtp_1 _166_ (.CLK(\CLKMUX.clk1 ),
    .D(_006_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\clk_div[5] ));
 sky130_fd_sc_hs__dfxtp_1 _167_ (.CLK(\CLKMUX.clk1 ),
    .D(_007_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\clk_div[6] ));
 sky130_fd_sc_hs__dfxtp_1 _168_ (.CLK(\CLKMUX.clk1 ),
    .D(_008_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\clk_div[7] ));
 sky130_fd_sc_hs__dfxtp_1 _169_ (.CLK(\CLKMUX.clk1 ),
    .D(_009_),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\clk_div[8] ));
 sky130_fd_sc_hs__dfxtp_1 _170_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[1] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[0] ));
 sky130_fd_sc_hs__dfxtp_1 _171_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[2] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[1] ));
 sky130_fd_sc_hs__dfxtp_1 _172_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[3] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[2] ));
 sky130_fd_sc_hs__dfxtp_1 _173_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[4] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[3] ));
 sky130_fd_sc_hs__dfxtp_1 _174_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[5] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[4] ));
 sky130_fd_sc_hs__dfxtp_1 _175_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[6] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[5] ));
 sky130_fd_sc_hs__dfxtp_1 _176_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[7] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[6] ));
 sky130_fd_sc_hs__dfxtp_1 _177_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[7] ));
 sky130_fd_sc_hs__dfxtp_1 _178_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[9] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[8] ));
 sky130_fd_sc_hs__dfxtp_1 _179_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[10] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[9] ));
 sky130_fd_sc_hs__dfxtp_1 _180_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[10] ));
 sky130_fd_sc_hs__dfxtp_1 _181_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[11] ));
 sky130_fd_sc_hs__dfxtp_1 _182_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[13] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[12] ));
 sky130_fd_sc_hs__dfxtp_1 _183_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[14] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[13] ));
 sky130_fd_sc_hs__dfxtp_1 _184_ (.CLK(\clk_div[8] ),
    .D(\shift_reg3[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[14] ));
 sky130_fd_sc_hs__dfxtp_1 _185_ (.CLK(\clk_div[8] ),
    .D(zero),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg3[15] ));
 sky130_fd_sc_hs__dfxtp_1 _186_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[1] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[0] ));
 sky130_fd_sc_hs__dfxtp_1 _187_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[2] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[1] ));
 sky130_fd_sc_hs__dfxtp_1 _188_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[3] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[2] ));
 sky130_fd_sc_hs__dfxtp_1 _189_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[4] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[3] ));
 sky130_fd_sc_hs__dfxtp_1 _190_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[5] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[4] ));
 sky130_fd_sc_hs__dfxtp_1 _191_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[6] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[5] ));
 sky130_fd_sc_hs__dfxtp_1 _192_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[7] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[6] ));
 sky130_fd_sc_hs__dfxtp_1 _193_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[7] ));
 sky130_fd_sc_hs__dfxtp_1 _194_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[9] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[8] ));
 sky130_fd_sc_hs__dfxtp_1 _195_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[10] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[9] ));
 sky130_fd_sc_hs__dfxtp_1 _196_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[10] ));
 sky130_fd_sc_hs__dfxtp_1 _197_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[11] ));
 sky130_fd_sc_hs__dfxtp_1 _198_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[13] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[12] ));
 sky130_fd_sc_hs__dfxtp_1 _199_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[14] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[13] ));
 sky130_fd_sc_hs__dfxtp_1 _200_ (.CLK(\clk_div[8] ),
    .D(\shift_reg2[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[14] ));
 sky130_fd_sc_hs__dfxtp_1 _201_ (.CLK(\clk_div[8] ),
    .D(one),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg2[15] ));
 sky130_fd_sc_hs__dfxtp_1 _202_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[1] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[0] ));
 sky130_fd_sc_hs__dfxtp_1 _203_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[2] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[1] ));
 sky130_fd_sc_hs__dfxtp_1 _204_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[3] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[2] ));
 sky130_fd_sc_hs__dfxtp_1 _205_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[4] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[3] ));
 sky130_fd_sc_hs__dfxtp_1 _206_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[5] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[4] ));
 sky130_fd_sc_hs__dfxtp_1 _207_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[6] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[5] ));
 sky130_fd_sc_hs__dfxtp_1 _208_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[7] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[6] ));
 sky130_fd_sc_hs__dfxtp_1 _209_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[7] ));
 sky130_fd_sc_hs__dfxtp_1 _210_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[9] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[8] ));
 sky130_fd_sc_hs__dfxtp_1 _211_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[10] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[9] ));
 sky130_fd_sc_hs__dfxtp_1 _212_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[10] ));
 sky130_fd_sc_hs__dfxtp_1 _213_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[11] ));
 sky130_fd_sc_hs__dfxtp_1 _214_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[13] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[12] ));
 sky130_fd_sc_hs__dfxtp_1 _215_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[14] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[13] ));
 sky130_fd_sc_hs__dfxtp_1 _216_ (.CLK(\clk_div[8] ),
    .D(\shift_reg1[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[14] ));
 sky130_fd_sc_hs__dfxtp_1 _217_ (.CLK(\clk_div[8] ),
    .D(zero),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg1[15] ));
 sky130_fd_sc_hs__dfxtp_1 _218_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[1] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[0] ));
 sky130_fd_sc_hs__dfxtp_1 _219_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[2] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[1] ));
 sky130_fd_sc_hs__dfxtp_1 _220_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[3] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[2] ));
 sky130_fd_sc_hs__dfxtp_1 _221_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[4] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[3] ));
 sky130_fd_sc_hs__dfxtp_1 _222_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[5] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[4] ));
 sky130_fd_sc_hs__dfxtp_1 _223_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[6] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[5] ));
 sky130_fd_sc_hs__dfxtp_1 _224_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[7] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[6] ));
 sky130_fd_sc_hs__dfxtp_1 _225_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[8] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[7] ));
 sky130_fd_sc_hs__dfxtp_1 _226_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[9] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[8] ));
 sky130_fd_sc_hs__dfxtp_1 _227_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[10] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[9] ));
 sky130_fd_sc_hs__dfxtp_1 _228_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[11] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[10] ));
 sky130_fd_sc_hs__dfxtp_1 _229_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[12] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[11] ));
 sky130_fd_sc_hs__dfxtp_1 _230_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[13] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[12] ));
 sky130_fd_sc_hs__dfxtp_1 _231_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[14] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[13] ));
 sky130_fd_sc_hs__dfxtp_1 _232_ (.CLK(\clk_div[8] ),
    .D(\shift_reg0[15] ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[14] ));
 sky130_fd_sc_hs__dfxtp_1 _233_ (.CLK(\clk_div[8] ),
    .D(one),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\shift_reg0[15] ));
 sky130_fd_sc_hs__dfrtp_1 _234_ (.CLK(_000_),
    .D(\CLKMUX.m3.Q2a ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m3.Q2b ));
 sky130_fd_sc_hs__dfrtn_1 _235_ (.CLK_N(_000_),
    .D(\CLKMUX.m3.q2a_in ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m3.Q2a ));
 sky130_fd_sc_hs__dfrtp_1 _236_ (.CLK(_001_),
    .D(\CLKMUX.m3.Q1a ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m3.Q1b ));
 sky130_fd_sc_hs__dfrtn_1 _237_ (.CLK_N(_001_),
    .D(\CLKMUX.m3.q1a_in ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m3.Q1a ));
 sky130_fd_sc_hs__dfrtn_1 _238_ (.CLK_N(\CLKMUX.clk4 ),
    .D(\CLKMUX.m2.Q2a ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m2.Q2b ));
 sky130_fd_sc_hs__dfrtp_1 _239_ (.CLK(\CLKMUX.clk4 ),
    .D(\CLKMUX.m2.q2a_in ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m2.Q2a ));
 sky130_fd_sc_hs__dfrtn_1 _240_ (.CLK_N(\CLKMUX.clk3 ),
    .D(\CLKMUX.m2.Q1a ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m2.Q1b ));
 sky130_fd_sc_hs__dfrtp_1 _241_ (.CLK(\CLKMUX.clk3 ),
    .D(\CLKMUX.m2.q1a_in ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m2.Q1a ));
 sky130_fd_sc_hs__dfrtn_1 _242_ (.CLK_N(\CLKMUX.clk2 ),
    .D(\CLKMUX.m1.Q2a ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m1.Q2b ));
 sky130_fd_sc_hs__dfrtp_1 _243_ (.CLK(\CLKMUX.clk2 ),
    .D(\CLKMUX.m1.q2a_in ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m1.Q2a ));
 sky130_fd_sc_hs__dfrtn_1 _244_ (.CLK_N(\CLKMUX.clk1 ),
    .D(\CLKMUX.m1.Q1a ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m1.Q1b ));
 sky130_fd_sc_hs__dfrtp_1 _245_ (.CLK(\CLKMUX.clk1 ),
    .D(\CLKMUX.m1.q1a_in ),
    .RESET_B(rst_n),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .Q(\CLKMUX.m1.Q1a ));
 sky130_fd_sc_hs__buf_2 _246_ (.A(\CLKMUX.clk2 ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(\clk_div[1] ));
 sky130_fd_sc_hs__buf_2 _247_ (.A(\CLKMUX.clk3 ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(\clk_div[2] ));
 sky130_fd_sc_hs__buf_2 _248_ (.A(\CLKMUX.clk4 ),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(\clk_div[3] ));
 sky130_fd_sc_hs__buf_2 _249_ (.A(clk_8mhz),
    .VGND(VGND),
  
    .VPWR(VPWR),
    .X(\clk_div[4] ));
 sky130_fd_sc_hs__decap_4 PHY_0 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_1 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_2 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_3 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_5 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_6 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_7 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_8 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_9 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_10 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_11 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_12 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_13 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_14 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_15 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_16 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_17 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_18 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_19 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_20 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_21 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_22 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_23 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_24 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_26 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_27 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_29 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_30 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_31 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_32 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_33 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_34 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_35 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_73 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_74 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_75 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_76 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_77 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_47 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_51 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_53 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_59 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_61 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_101 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_105 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_107 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_113 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_115 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_133 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_155 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_159 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_161 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_171 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_179 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_187 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_198 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_206 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_214 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_1_6 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_24 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_45 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_52 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_63 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_1_67 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_85 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_106 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_113 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_1_115 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_133 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_160 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_170 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_174 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_199 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_207 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_47 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_58 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_101 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_2_105 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_112 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_133 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_155 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_2_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_187 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_198 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_205 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_213 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_29 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_50 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_3_59 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_66 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_76 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_97 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_106 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_117 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_124 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_145 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_156 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_160 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_3_167 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_171 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_3_179 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_203 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_210 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_3_214 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_36 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_40 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_4_42 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_60 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_69 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_101 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_110 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_121 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_125 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_133 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_4_155 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_4_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_187 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_197 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_4_204 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_212 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_4_214 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_10 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_31 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_52 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_63 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_67 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_76 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_97 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_105 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_5_107 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_128 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_132 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_140 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_148 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_155 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_159 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_5_161 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_5_165 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_189 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_5_193 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_5_205 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_213 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_38 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_59 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_69 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_73 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_75 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_86 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_95 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_99 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_107 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_128 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_132 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_134 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_144 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_148 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_172 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_182 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_186 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_188 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_6_205 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_213 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_8 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_10 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_17 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_38 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_42 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_50 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_62 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_7_69 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_77 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_81 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_86 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_95 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_106 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_113 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_131 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_152 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_159 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_161 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_170 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_174 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_198 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_213 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_8_30 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_37 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_41 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_49 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_8_57 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_65 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_75 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_8_101 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_8_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_8_127 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_145 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_154 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_8_181 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_8_205 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_213 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_9_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_9_12 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_20 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_24 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_9_26 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_44 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_52 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_9_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_63 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_9_67 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_85 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_106 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_9_113 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_9_122 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_130 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_149 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_159 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_9_161 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_188 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_192 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_9_205 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_213 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_10_30 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_37 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_58 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_86 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_10_88 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_106 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_10_116 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_124 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_133 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_10_145 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_10_153 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_177 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_187 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_10_205 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_213 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_11_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_29 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_50 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_11_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_64 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_74 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_85 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_11_106 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_11_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_11_117 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_128 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_149 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_158 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_11_167 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_192 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_11_207 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_47 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_57 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_12_64 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_72 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_12_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_107 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_12_114 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_122 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_12_124 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_128 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_132 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_12_134 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_155 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_162 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_12_166 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_12_172 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_12_180 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_12_188 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_12_205 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_213 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_12 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_20 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_24 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_43 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_52 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_63 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_13_65 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_83 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_104 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_117 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_138 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_147 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_155 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_159 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_13_161 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_168 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_176 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_184 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_188 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_13_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_197 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_205 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_213 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_49 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_58 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_92 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_102 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_110 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_114 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_133 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_145 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_153 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_161 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_169 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_177 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_185 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_198 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_206 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_14_214 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_15_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_15_6 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_15_10 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_15_31 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_15_52 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_15_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_15_59 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_15_78 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_15_99 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_15_106 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_15_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_15_117 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_15_138 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_15_147 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_15_155 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_15_159 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_15_161 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_15_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_15_171 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_15_179 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_15_187 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_15_195 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_15_203 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_15_211 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_16_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_16_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_16_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_16_47 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_16_51 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_16_53 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_16_58 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_16_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_16_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_91 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_16_99 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_16_117 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_16_121 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_16_129 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_16_133 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_144 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_152 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_160 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_168 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_176 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_16_184 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_16_188 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_198 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_16_206 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_16_214 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_4 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_12 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_17_25 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_17_28 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_17_37 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_17_47 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_17_51 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_17_53 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_17_55 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_17_57 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_17_75 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_17_79 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_17_82 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_17_91 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_99 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_17_107 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_109 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_117 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_125 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_17_133 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_136 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_144 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_152 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_17_160 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_163 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_171 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_179 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_17_187 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_190 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_198 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_17_206 (.VGND(VGND),
  
    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_17_214 (.VGND(VGND),
  
    .VPWR(VPWR));
endmodule
