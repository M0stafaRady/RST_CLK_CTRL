module freq_mul_x8 (clk_out,
    clk_ref,
    en,
    fb_in,
    fb_out,
    rst_n,
    VGND,
    VPWR,
    trim);
 output clk_out;
 input clk_ref;
 input en;
 input fb_in;
 output fb_out;
 input rst_n;
 input VGND;
 input VPWR;
 input [1:0] trim;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire \clk_out_half_cntr[0] ;
 wire \clk_out_half_cntr[1] ;
 wire \clk_out_half_cntr[2] ;
 wire \clk_out_half_cntr[3] ;
 wire \clk_out_half_width[0] ;
 wire \clk_out_half_width[1] ;
 wire \clk_out_half_width[2] ;
 wire \clk_out_half_width[3] ;
 wire \clk_out_half_width[4] ;
 wire \clk_out_half_width[5] ;
 wire \clk_out_half_width_rem[1] ;
 wire \clk_out_half_width_rem[2] ;
 wire \clk_out_half_width_rem[3] ;
 wire clk_ref_sync;
 wire clk_ref_sync_dly;
 wire \clk_ref_sync_ff[0] ;
 wire \clk_ref_sync_width[0] ;
 wire \clk_ref_sync_width[1] ;
 wire \clk_ref_sync_width[2] ;
 wire \clk_ref_sync_width[3] ;
 wire \clk_ref_sync_width[4] ;
 wire \clk_ref_sync_width[5] ;
 wire \clk_ref_sync_width[6] ;
 wire \clk_ref_sync_width[7] ;
 wire \clk_ref_sync_width[8] ;
 wire \clk_ref_sync_width[9] ;
 wire \half_cyc_cntr[0] ;
 wire \half_cyc_cntr[1] ;
 wire \half_cyc_cntr[2] ;
 wire \half_cyc_cntr[3] ;
 wire \half_cyc_cntr[4] ;
 wire \half_cyc_cntr[5] ;
 wire \rosc.chain_2[1] ;
 wire \rosc.chain_2[2] ;
 wire \rosc.chain_4[1] ;
 wire \rosc.chain_4[2] ;
 wire \rosc.chain_4[3] ;
 wire \rosc.chain_4[4] ;
 wire \rosc.chain_6[1] ;
 wire \rosc.chain_6[2] ;
 wire \rosc.chain_6[3] ;
 wire \rosc.chain_6[4] ;
 wire \rosc.chain_6[5] ;
 wire \rosc.chain_6[6] ;
 wire \rosc.clk ;
 wire \rosc.inv_out[0] ;
 wire \rosc.inv_out[1] ;
 wire \rosc.mux_out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;

 sky130_fd_sc_hs__nor2b_2 _070_ (.A(clk_ref_sync_dly),
    .B_N(clk_ref_sync),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_047_));
 sky130_fd_sc_hs__and2_1 _071_ (.A(\clk_out_half_cntr[2] ),
    .B(\clk_out_half_cntr[3] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_048_));
 sky130_fd_sc_hs__nand3_2 _072_ (.A(\clk_out_half_cntr[0] ),
    .B(\clk_out_half_cntr[1] ),
    .C(\clk_out_half_width_rem[1] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_049_));
 sky130_fd_sc_hs__nand2b_1 _073_ (.A_N(\clk_out_half_cntr[0] ),
    .B(\clk_out_half_width_rem[3] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_050_));
 sky130_fd_sc_hs__nand3b_1 _074_ (.A_N(\clk_out_half_cntr[1] ),
    .B(\clk_out_half_width_rem[2] ),
    .C(\clk_out_half_cntr[0] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_051_));
 sky130_fd_sc_hs__o211ai_4 _075_ (.A1(_048_),
    .A2(_049_),
    .B1(_050_),
    .C1(_051_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_052_));
 sky130_fd_sc_hs__nor2_1 _076_ (.A(\half_cyc_cntr[2] ),
    .B(\half_cyc_cntr[5] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_053_));
 sky130_fd_sc_hs__nor2_4 _077_ (.A(\half_cyc_cntr[3] ),
    .B(\half_cyc_cntr[4] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_054_));
 sky130_fd_sc_hs__nand4b_4 _078_ (.A_N(\half_cyc_cntr[1] ),
    .B(_053_),
    .C(_054_),
    .D(\half_cyc_cntr[0] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_055_));
 sky130_fd_sc_hs__nor3_4 _079_ (.A(\half_cyc_cntr[0] ),
    .B(\half_cyc_cntr[1] ),
    .C(\half_cyc_cntr[2] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_056_));
 sky130_fd_sc_hs__nand2_1 _080_ (.A(_054_),
    .B(_056_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_057_));
 sky130_fd_sc_hs__nand3b_2 _081_ (.A_N(\half_cyc_cntr[5] ),
    .B(_054_),
    .C(_056_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_058_));
 sky130_fd_sc_hs__mux2i_4 _082_ (.A0(_055_),
    .A1(_058_),
    .S(_052_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_059_));
 sky130_fd_sc_hs__nor2_4 _083_ (.A(net10),
    .B(_059_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_060_));
 sky130_fd_sc_hs__o21ai_1 _084_ (.A1(net10),
    .A2(_059_),
    .B1(\clk_out_half_width[0] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_061_));
 sky130_fd_sc_hs__o31ai_1 _085_ (.A1(\half_cyc_cntr[0] ),
    .A2(net10),
    .A3(_059_),
    .B1(_061_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_000_));
 sky130_fd_sc_hs__xnor2_1 _086_ (.A(\half_cyc_cntr[0] ),
    .B(\half_cyc_cntr[1] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_062_));
 sky130_fd_sc_hs__mux2_1 _087_ (.A0(\clk_out_half_width[1] ),
    .A1(_062_),
    .S(_060_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_001_));
 sky130_fd_sc_hs__o21ai_1 _088_ (.A1(\half_cyc_cntr[0] ),
    .A2(\half_cyc_cntr[1] ),
    .B1(\half_cyc_cntr[2] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_063_));
 sky130_fd_sc_hs__nand2b_1 _089_ (.A_N(_056_),
    .B(_063_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_064_));
 sky130_fd_sc_hs__mux2_1 _090_ (.A0(\clk_out_half_width[2] ),
    .A1(_064_),
    .S(_060_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_002_));
 sky130_fd_sc_hs__xor2_1 _091_ (.A(\half_cyc_cntr[3] ),
    .B(_056_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_065_));
 sky130_fd_sc_hs__mux2_1 _092_ (.A0(\clk_out_half_width[3] ),
    .A1(_065_),
    .S(_060_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_003_));
 sky130_fd_sc_hs__o41ai_1 _093_ (.A1(\half_cyc_cntr[0] ),
    .A2(\half_cyc_cntr[1] ),
    .A3(\half_cyc_cntr[3] ),
    .A4(\half_cyc_cntr[2] ),
    .B1(\half_cyc_cntr[4] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_066_));
 sky130_fd_sc_hs__nand2_1 _094_ (.A(_057_),
    .B(_066_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_067_));
 sky130_fd_sc_hs__mux2_1 _095_ (.A0(\clk_out_half_width[4] ),
    .A1(_067_),
    .S(_060_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_004_));
 sky130_fd_sc_hs__nand2_1 _096_ (.A(\half_cyc_cntr[5] ),
    .B(_057_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_068_));
 sky130_fd_sc_hs__nand2_1 _097_ (.A(_058_),
    .B(_068_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_069_));
 sky130_fd_sc_hs__mux2_1 _098_ (.A0(\clk_out_half_width[5] ),
    .A1(_069_),
    .S(_060_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hs__mux2_1 _099_ (.A0(\clk_out_half_width_rem[1] ),
    .A1(\clk_ref_sync_width[1] ),
    .S(net9),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hs__mux2_1 _100_ (.A0(\clk_out_half_width_rem[2] ),
    .A1(\clk_ref_sync_width[2] ),
    .S(net9),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_007_));
 sky130_fd_sc_hs__mux2_1 _101_ (.A0(\clk_out_half_width_rem[3] ),
    .A1(\clk_ref_sync_width[3] ),
    .S(net9),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_008_));
 sky130_fd_sc_hs__mux2_1 _102_ (.A0(\clk_out_half_width[0] ),
    .A1(\clk_ref_sync_width[4] ),
    .S(net10),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_009_));
 sky130_fd_sc_hs__mux2_1 _103_ (.A0(\clk_out_half_width[1] ),
    .A1(\clk_ref_sync_width[5] ),
    .S(net10),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_010_));
 sky130_fd_sc_hs__mux2_1 _104_ (.A0(\clk_out_half_width[2] ),
    .A1(\clk_ref_sync_width[6] ),
    .S(net10),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_011_));
 sky130_fd_sc_hs__mux2_1 _105_ (.A0(\clk_out_half_width[3] ),
    .A1(\clk_ref_sync_width[7] ),
    .S(net10),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_012_));
 sky130_fd_sc_hs__mux2_1 _106_ (.A0(\clk_out_half_width[4] ),
    .A1(\clk_ref_sync_width[8] ),
    .S(net10),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_013_));
 sky130_fd_sc_hs__mux2_1 _107_ (.A0(\clk_out_half_width[5] ),
    .A1(\clk_ref_sync_width[9] ),
    .S(_047_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hs__nand2_1 _108_ (.A(\clk_out_half_cntr[0] ),
    .B(_059_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_030_));
 sky130_fd_sc_hs__xor2_1 _109_ (.A(\clk_out_half_cntr[0] ),
    .B(_059_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_015_));
 sky130_fd_sc_hs__xnor2_1 _110_ (.A(\clk_out_half_cntr[1] ),
    .B(_030_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_016_));
 sky130_fd_sc_hs__a31oi_1 _111_ (.A1(\clk_out_half_cntr[0] ),
    .A2(\clk_out_half_cntr[1] ),
    .A3(_059_),
    .B1(\clk_out_half_cntr[2] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_031_));
 sky130_fd_sc_hs__nand4_2 _112_ (.A(\clk_out_half_cntr[0] ),
    .B(\clk_out_half_cntr[1] ),
    .C(\clk_out_half_cntr[2] ),
    .D(_059_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_032_));
 sky130_fd_sc_hs__nor2b_1 _113_ (.A(_031_),
    .B_N(_032_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_017_));
 sky130_fd_sc_hs__xnor2_1 _114_ (.A(\clk_out_half_cntr[3] ),
    .B(_032_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_018_));
 sky130_fd_sc_hs__xor2_1 _115_ (.A(net7),
    .B(_059_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_019_));
 sky130_fd_sc_hs__nor2_1 _116_ (.A(\clk_ref_sync_width[0] ),
    .B(net9),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_020_));
 sky130_fd_sc_hs__a21oi_1 _117_ (.A1(\clk_ref_sync_width[0] ),
    .A2(\clk_ref_sync_width[1] ),
    .B1(net9),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_033_));
 sky130_fd_sc_hs__o21a_1 _118_ (.A1(\clk_ref_sync_width[0] ),
    .A2(\clk_ref_sync_width[1] ),
    .B1(_033_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_021_));
 sky130_fd_sc_hs__a21oi_1 _119_ (.A1(\clk_ref_sync_width[0] ),
    .A2(\clk_ref_sync_width[1] ),
    .B1(\clk_ref_sync_width[2] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_034_));
 sky130_fd_sc_hs__and3_1 _120_ (.A(\clk_ref_sync_width[0] ),
    .B(\clk_ref_sync_width[1] ),
    .C(\clk_ref_sync_width[2] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_035_));
 sky130_fd_sc_hs__nor3_1 _121_ (.A(net9),
    .B(_034_),
    .C(_035_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_022_));
 sky130_fd_sc_hs__nor2_1 _122_ (.A(\clk_ref_sync_width[3] ),
    .B(_035_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_036_));
 sky130_fd_sc_hs__and4_1 _123_ (.A(\clk_ref_sync_width[0] ),
    .B(\clk_ref_sync_width[1] ),
    .C(\clk_ref_sync_width[2] ),
    .D(\clk_ref_sync_width[3] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_037_));
 sky130_fd_sc_hs__nor3_1 _124_ (.A(net9),
    .B(_036_),
    .C(_037_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_023_));
 sky130_fd_sc_hs__a21oi_1 _125_ (.A1(\clk_ref_sync_width[4] ),
    .A2(_037_),
    .B1(net9),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_038_));
 sky130_fd_sc_hs__o21a_1 _126_ (.A1(\clk_ref_sync_width[4] ),
    .A2(_037_),
    .B1(_038_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_024_));
 sky130_fd_sc_hs__a21oi_1 _127_ (.A1(\clk_ref_sync_width[4] ),
    .A2(_037_),
    .B1(\clk_ref_sync_width[5] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_039_));
 sky130_fd_sc_hs__and3_1 _128_ (.A(\clk_ref_sync_width[4] ),
    .B(\clk_ref_sync_width[5] ),
    .C(_037_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_040_));
 sky130_fd_sc_hs__nor3_1 _129_ (.A(net9),
    .B(_039_),
    .C(_040_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_025_));
 sky130_fd_sc_hs__a21oi_1 _130_ (.A1(\clk_ref_sync_width[6] ),
    .A2(_040_),
    .B1(net9),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_041_));
 sky130_fd_sc_hs__o21a_1 _131_ (.A1(\clk_ref_sync_width[6] ),
    .A2(_040_),
    .B1(_041_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_026_));
 sky130_fd_sc_hs__a21oi_1 _132_ (.A1(\clk_ref_sync_width[6] ),
    .A2(_040_),
    .B1(\clk_ref_sync_width[7] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_042_));
 sky130_fd_sc_hs__and3_1 _133_ (.A(\clk_ref_sync_width[6] ),
    .B(\clk_ref_sync_width[7] ),
    .C(_040_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_043_));
 sky130_fd_sc_hs__nor3_1 _134_ (.A(_047_),
    .B(_042_),
    .C(_043_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_027_));
 sky130_fd_sc_hs__a21oi_1 _135_ (.A1(\clk_ref_sync_width[8] ),
    .A2(_043_),
    .B1(net10),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_044_));
 sky130_fd_sc_hs__o21a_1 _136_ (.A1(\clk_ref_sync_width[8] ),
    .A2(_043_),
    .B1(_044_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_028_));
 sky130_fd_sc_hs__a21oi_1 _137_ (.A1(\clk_ref_sync_width[8] ),
    .A2(_043_),
    .B1(\clk_ref_sync_width[9] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_045_));
 sky130_fd_sc_hs__and3_1 _138_ (.A(\clk_ref_sync_width[8] ),
    .B(\clk_ref_sync_width[9] ),
    .C(_043_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(_046_));
 sky130_fd_sc_hs__nor3_1 _139_ (.A(_047_),
    .B(_045_),
    .C(_046_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(_029_));
 sky130_fd_sc_hs__dfxtp_1 _140_ (.CLK(net13),
    .D(net1),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_ff[0] ));
 sky130_fd_sc_hs__dfxtp_1 _141_ (.CLK(net13),
    .D(\clk_ref_sync_ff[0] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(clk_ref_sync));
 sky130_fd_sc_hs__dfxtp_1 _142_ (.CLK(net13),
    .D(clk_ref_sync),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(clk_ref_sync_dly));
 sky130_fd_sc_hs__dfxtp_1 _143_ (.CLK(net11),
    .D(_006_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_width_rem[1] ));
 sky130_fd_sc_hs__dfxtp_1 _144_ (.CLK(net11),
    .D(_007_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_width_rem[2] ));
 sky130_fd_sc_hs__dfxtp_1 _145_ (.CLK(net11),
    .D(_008_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_width_rem[3] ));
 sky130_fd_sc_hs__dfxtp_1 _146_ (.CLK(net11),
    .D(_009_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_width[0] ));
 sky130_fd_sc_hs__dfxtp_1 _147_ (.CLK(net12),
    .D(_010_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_width[1] ));
 sky130_fd_sc_hs__dfxtp_1 _148_ (.CLK(net13),
    .D(_011_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_width[2] ));
 sky130_fd_sc_hs__dfxtp_1 _149_ (.CLK(net13),
    .D(_012_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_width[3] ));
 sky130_fd_sc_hs__dfxtp_1 _150_ (.CLK(net13),
    .D(_013_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_width[4] ));
 sky130_fd_sc_hs__dfxtp_1 _151_ (.CLK(net13),
    .D(_014_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_width[5] ));
 sky130_fd_sc_hs__dfrtp_2 _152_ (.CLK(net13),
    .D(_015_),
    .RESET_B(net4),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_cntr[0] ));
 sky130_fd_sc_hs__dfrtp_2 _153_ (.CLK(net11),
    .D(_016_),
    .RESET_B(net4),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_cntr[1] ));
 sky130_fd_sc_hs__dfrtp_1 _154_ (.CLK(net12),
    .D(_017_),
    .RESET_B(net4),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_cntr[2] ));
 sky130_fd_sc_hs__dfrtp_1 _155_ (.CLK(net14),
    .D(_018_),
    .RESET_B(net4),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_out_half_cntr[3] ));
 sky130_fd_sc_hs__dfrtp_1 _156_ (.CLK(net14),
    .D(_019_),
    .RESET_B(net4),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(net7));
 sky130_fd_sc_hs__dfxtp_2 _157_ (.CLK(net14),
    .D(_000_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\half_cyc_cntr[0] ));
 sky130_fd_sc_hs__dfxtp_2 _158_ (.CLK(net14),
    .D(_001_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\half_cyc_cntr[1] ));
 sky130_fd_sc_hs__dfxtp_2 _159_ (.CLK(net14),
    .D(_002_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\half_cyc_cntr[2] ));
 sky130_fd_sc_hs__dfxtp_1 _160_ (.CLK(net14),
    .D(_003_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\half_cyc_cntr[3] ));
 sky130_fd_sc_hs__dfxtp_1 _161_ (.CLK(net14),
    .D(_004_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\half_cyc_cntr[4] ));
 sky130_fd_sc_hs__dfxtp_1 _162_ (.CLK(net14),
    .D(_005_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\half_cyc_cntr[5] ));
 sky130_fd_sc_hs__dfxtp_1 _163_ (.CLK(net12),
    .D(_020_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[0] ));
 sky130_fd_sc_hs__dfxtp_1 _164_ (.CLK(net11),
    .D(_021_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[1] ));
 sky130_fd_sc_hs__dfxtp_1 _165_ (.CLK(net11),
    .D(_022_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[2] ));
 sky130_fd_sc_hs__dfxtp_1 _166_ (.CLK(net11),
    .D(_023_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[3] ));
 sky130_fd_sc_hs__dfxtp_1 _167_ (.CLK(net11),
    .D(_024_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[4] ));
 sky130_fd_sc_hs__dfxtp_1 _168_ (.CLK(net11),
    .D(_025_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[5] ));
 sky130_fd_sc_hs__dfxtp_1 _169_ (.CLK(net12),
    .D(_026_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[6] ));
 sky130_fd_sc_hs__dfxtp_1 _170_ (.CLK(net12),
    .D(_027_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[7] ));
 sky130_fd_sc_hs__dfxtp_1 _171_ (.CLK(net13),
    .D(_028_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[8] ));
 sky130_fd_sc_hs__dfxtp_1 _172_ (.CLK(net13),
    .D(_029_),
    .VGND(VGND),

    .VPWR(VPWR),
    .Q(\clk_ref_sync_width[9] ));
 sky130_fd_sc_hs__dlymetal6s2s_1 \rosc.BUF  (.A(net8),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(\rosc.clk ));
 sky130_fd_sc_hs__nand2_2 \rosc.ENABLE  (.A(net2),
    .B(\rosc.inv_out[1] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(net8));
 sky130_fd_sc_hs__inv_2 \rosc.INV_0  (.A(\rosc.mux_out ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.inv_out[0] ));
 sky130_fd_sc_hs__inv_2 \rosc.INV_1  (.A(\rosc.inv_out[0] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.inv_out[1] ));
 sky130_fd_sc_hs__inv_1 \rosc.INV_CHAIN_2_0  (.A(net3),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_2[1] ));
 sky130_fd_sc_hs__inv_1 \rosc.INV_CHAIN_2_1  (.A(\rosc.chain_2[1] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_2[2] ));
 sky130_fd_sc_hs__inv_1 \rosc.INV_CHAIN_4_0  (.A(net3),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_4[1] ));
 sky130_fd_sc_hs__inv_1 \rosc.INV_CHAIN_4_1  (.A(\rosc.chain_4[1] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_4[2] ));
 sky130_fd_sc_hs__inv_1 \rosc.INV_CHAIN_4_2  (.A(\rosc.chain_4[2] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_4[3] ));
 sky130_fd_sc_hs__inv_1 \rosc.INV_CHAIN_4_3  (.A(\rosc.chain_4[3] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_4[4] ));
 sky130_fd_sc_hs__inv_4 \rosc.INV_CHAIN_6_0  (.A(net3),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_6[1] ));
 sky130_fd_sc_hs__inv_2 \rosc.INV_CHAIN_6_1  (.A(\rosc.chain_6[1] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_6[2] ));
 sky130_fd_sc_hs__inv_2 \rosc.INV_CHAIN_6_2  (.A(\rosc.chain_6[2] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_6[3] ));
 sky130_fd_sc_hs__inv_2 \rosc.INV_CHAIN_6_3  (.A(\rosc.chain_6[3] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_6[4] ));
 sky130_fd_sc_hs__inv_2 \rosc.INV_CHAIN_6_4  (.A(\rosc.chain_6[4] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_6[5] ));
 sky130_fd_sc_hs__inv_2 \rosc.INV_CHAIN_6_5  (.A(\rosc.chain_6[5] ),
    .VGND(VGND),

    .VPWR(VPWR),
    .Y(\rosc.chain_6[6] ));
 sky130_fd_sc_hs__mux4_1 \rosc.MUX  (.A0(net3),
    .A1(\rosc.chain_2[2] ),
    .A2(\rosc.chain_4[4] ),
    .A3(\rosc.chain_6[6] ),
    .S0(net5),
    .S1(net6),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(\rosc.mux_out ));
 sky130_fd_sc_hs__decap_4 PHY_0 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_1 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_2 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_3 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_5 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_6 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_7 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_8 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_9 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_10 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_11 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_13 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_14 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_15 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_16 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_17 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_18 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_19 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_20 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_21 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_22 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_23 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_24 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_25 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_26 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_27 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 PHY_29 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_30 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_31 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_32 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_33 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_34 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_35 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_36 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_37 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_38 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_39 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_40 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_41 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_42 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_43 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_44 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_45 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_46 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_47 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_48 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_49 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_50 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_51 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_52 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_53 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_54 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_55 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_56 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_57 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_58 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_59 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_60 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_61 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_62 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_63 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_64 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_65 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_66 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_67 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_68 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_69 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_70 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_71 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_72 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_73 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_74 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_75 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_76 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_77 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hs__clkbuf_1 input1 (.A(clk_ref),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hs__clkbuf_1 input2 (.A(en),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hs__buf_8 input3 (.A(fb_in),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hs__clkbuf_4 input4 (.A(rst_n),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hs__clkbuf_1 input5 (.A(trim[0]),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hs__clkbuf_1 input6 (.A(trim[1]),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hs__buf_4 output7 (.A(net7),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(clk_out));
 sky130_fd_sc_hs__buf_8 output8 (.A(net8),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(fb_out));
 sky130_fd_sc_hs__clkbuf_4 fanout9 (.A(net10),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hs__buf_4 fanout10 (.A(_047_),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hs__clkbuf_4 fanout11 (.A(net12),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hs__buf_2 fanout12 (.A(\rosc.clk ),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hs__clkbuf_4 fanout13 (.A(\rosc.clk ),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hs__buf_2 fanout14 (.A(\rosc.clk ),
    .VGND(VGND),

    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hs__fill_8 FILLER_0_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_16 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_21 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_25 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_36 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_44 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_52 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_0_55 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_63 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_69 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_73 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_75 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_79 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_82 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_86 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_91 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_98 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_105 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_107 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_109 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_117 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_121 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_133 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_136 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_140 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_159 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_161 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_0_163 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_0_169 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_0_173 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_20 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_36 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_44 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_52 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_55 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_63 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_71 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_1_79 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_83 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_90 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_99 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_106 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_109 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_114 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_1_121 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_125 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_133 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_141 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_160 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_1_163 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_1_171 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_1_173 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_20 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_24 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_2_26 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_36 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_44 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_52 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_60 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_68 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_76 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_2_80 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_82 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_93 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_117 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_125 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_2_133 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_2_136 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_161 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_2_169 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_2_173 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_20 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_36 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_44 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_52 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_55 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_63 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_69 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_77 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_84 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_3_92 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_100 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_105 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_3_107 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_109 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_116 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_137 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_3_144 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_160 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_163 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_3_172 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_4_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_4_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_20 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_24 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_4_26 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_4_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_4_36 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_4_44 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_4_52 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_60 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_4_64 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_69 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_79 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_82 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_4_86 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_93 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_114 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_121 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_4_125 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_133 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_136 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_147 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_4_168 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_4_172 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_5_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_5_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_5_20 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_5_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_5_36 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_5_44 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_52 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_55 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_5_59 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_77 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_98 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_106 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_109 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_120 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_5_124 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_131 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_152 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_160 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_5_163 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_5_169 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_5_173 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_6_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_6_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_20 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_25 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_34 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_6_41 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_49 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_54 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_6_63 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_71 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_77 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_82 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_90 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_6_111 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_119 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_121 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_130 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_134 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_136 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_141 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_6_162 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_6_171 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_6_173 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_8 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_33 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_7_41 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_49 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_53 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_7_55 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_63 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_7_81 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_89 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_91 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_101 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_105 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_107 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_109 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_111 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_129 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_133 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_143 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_7_156 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_160 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_7_163 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_7_171 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_7_173 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_25 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_47 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_8_51 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_58 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_79 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_82 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_8_90 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_8_98 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_108 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_130 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_8_134 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_136 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_147 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_8_168 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_8_172 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_9_6 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_13 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_34 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_38 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_9_40 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_50 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_55 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_63 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_9_67 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_74 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_78 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_97 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_106 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_109 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_120 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_124 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_9_126 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_145 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_9_158 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_163 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_9_172 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_8 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_10_10 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_15 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_25 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_10_30 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_38 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_59 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_66 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_79 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_82 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_101 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_110 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_114 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_133 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_136 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_10_157 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_161 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_10_172 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_11_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_11_16 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_34 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_47 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_11_51 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_11_53 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_11_55 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_86 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_99 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_11_106 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_109 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_11_113 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_128 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_153 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_11_160 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_11_163 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_11_170 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_25 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_39 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_43 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_12_52 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_60 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_79 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_82 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_89 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_116 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_129 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_133 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_136 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_12_156 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_12_172 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_16 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_24 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_52 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_55 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_62 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_74 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_102 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_106 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_109 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_13_117 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_127 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_13_154 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_163 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_13_168 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_13_172 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_4 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_12 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_16 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_14_18 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_25 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_28 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_36 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_45 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_14_53 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_55 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_14_63 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_74 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_78 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_14_80 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_82 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_91 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_14_99 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_106 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_109 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_117 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_14_119 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_8 FILLER_14_127 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_136 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_146 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_157 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_1 FILLER_14_161 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_163 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__decap_4 FILLER_14_168 (.VGND(VGND),

    .VPWR(VPWR));
 sky130_fd_sc_hs__fill_2 FILLER_14_172 (.VGND(VGND),

    .VPWR(VPWR));
endmodule
